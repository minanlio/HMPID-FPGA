-- megafunction wizard: %ALTREMOTE_UPDATE%CBX%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altremote_update 

-- ============================================================
-- File Name: alt_remote.vhd
-- Megafunction Name(s):
-- 			altremote_update
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 6.0 Build 202 06/20/2006 SP 1 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2006 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--altremote_update DEVICE_FAMILY="Stratix II" operation_mode="local" sim_init_config="application" sim_init_page_select=1 sim_init_status=15 busy clock data_out param pgmout read_param reconfig reset reset_timer
--VERSION_BEGIN 6.0 cbx_altremote_update 2005:11:22:18:11:24:SJ cbx_cycloneii 2006:02:07:15:19:20:SJ cbx_lpm_add_sub 2006:01:09:11:17:20:SJ cbx_lpm_compare 2006:01:09:11:15:40:SJ cbx_lpm_counter 2006:03:23:14:19:24:SJ cbx_lpm_decode 2006:01:09:11:16:44:SJ cbx_mgl 2006:05:17:10:06:16:SJ cbx_stratix 2006:05:17:09:28:32:SJ cbx_stratixii 2006:03:03:09:35:36:SJ  VERSION_END


--lpm_counter DEVICE_FAMILY="Stratix II" lpm_direction="UP" lpm_width=5 clock cnt_en q sclr
--VERSION_BEGIN 6.0 cbx_cycloneii 2006:02:07:15:19:20:SJ cbx_lpm_add_sub 2006:01:09:11:17:20:SJ cbx_lpm_compare 2006:01:09:11:15:40:SJ cbx_lpm_counter 2006:03:23:14:19:24:SJ cbx_lpm_decode 2006:01:09:11:16:44:SJ cbx_mgl 2006:05:17:10:06:16:SJ cbx_stratix 2006:05:17:09:28:32:SJ cbx_stratixii 2006:03:03:09:35:36:SJ  VERSION_END

 LIBRARY stratixii;
 USE stratixii.all;

--synthesis_resources = lut 5 reg 5 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  alt_remote_cntr_c88 IS 
	 PORT 
	 ( 
		 clock	:	IN  STD_LOGIC;
		 cnt_en	:	IN  STD_LOGIC := '1';
		 q	:	OUT  STD_LOGIC_VECTOR (4 DOWNTO 0);
		 sclr	:	IN  STD_LOGIC := '0'
	 ); 
 END alt_remote_cntr_c88;

 ARCHITECTURE RTL OF alt_remote_cntr_c88 IS

	 ATTRIBUTE synthesis_clearbox : boolean;
	 ATTRIBUTE synthesis_clearbox OF RTL : ARCHITECTURE IS true;
	 SIGNAL  wire_counter_comb_bita_0cout	:	STD_LOGIC;
	 SIGNAL  wire_counter_comb_bita_1cout	:	STD_LOGIC;
	 SIGNAL  wire_counter_comb_bita_2cout	:	STD_LOGIC;
	 SIGNAL  wire_counter_comb_bita_3cout	:	STD_LOGIC;
	 SIGNAL  wire_counter_comb_bita_0sumout	:	STD_LOGIC;
	 SIGNAL  wire_counter_comb_bita_1sumout	:	STD_LOGIC;
	 SIGNAL  wire_counter_comb_bita_2sumout	:	STD_LOGIC;
	 SIGNAL  wire_counter_comb_bita_3sumout	:	STD_LOGIC;
	 SIGNAL  wire_counter_comb_bita_4sumout	:	STD_LOGIC;
	 SIGNAL  wire_counter_reg_bit20a_adatasdata	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_counter_reg_bit20a_ena	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_counter_reg_bit20a_regout	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_counter_reg_bit20a_sload	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_cntr2_w_lg_w_lg_sset334w335w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_cntr2_w_lg_clk_en342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cntr2_w_lg_sset336w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_cntr2_w_lg_external_cin332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cntr2_w_lg_sset334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cntr2_w_lg_w_lg_sset336w337w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_cntr2_w_lg_w_lg_w_lg_cnt_en339w340w341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cntr2_w_lg_w_lg_cnt_en339w340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cntr2_w_lg_cnt_en339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cntr2_w_lg_sset338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  aclr_actual :	STD_LOGIC;
	 SIGNAL  clk_en	:	STD_LOGIC;
	 SIGNAL  data	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  external_cin :	STD_LOGIC;
	 SIGNAL  lsb_cin :	STD_LOGIC;
	 SIGNAL  s_val :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  safe_q :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  sload	:	STD_LOGIC;
	 SIGNAL  sset	:	STD_LOGIC;
	 SIGNAL  updown_dir :	STD_LOGIC;
	 SIGNAL  updown_lsb :	STD_LOGIC;
	 SIGNAL  updown_other_bits :	STD_LOGIC;
	 COMPONENT  stratixii_lcell_comb
	 GENERIC 
	 (
		EXTENDED_LUT	:	STRING := "OFF";
		LUT_MASK	:	STD_LOGIC_VECTOR(63 DOWNTO 0);
		SHARED_ARITH	:	STRING := "OFF";
		lpm_type	:	STRING := "stratixii_lcell_comb"
	 );
	 PORT
	 ( 
		cin	:	IN STD_LOGIC := '0';
		combout	:	OUT STD_LOGIC;
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC := '0';
		datab	:	IN STD_LOGIC := '0';
		datac	:	IN STD_LOGIC := '0';
		datad	:	IN STD_LOGIC := '0';
		datae	:	IN STD_LOGIC := '0';
		dataf	:	IN STD_LOGIC := '0';
		datag	:	IN STD_LOGIC := '0';
		sharein	:	IN STD_LOGIC := '0';
		shareout	:	OUT STD_LOGIC;
		sumout	:	OUT STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  stratixii_lcell_ff
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		adatasdata	:	IN STD_LOGIC := '0';
		aload	:	IN STD_LOGIC := '0';
		clk	:	IN STD_LOGIC;
		datain	:	IN STD_LOGIC;
		ena	:	IN STD_LOGIC := '1';
		regout	:	OUT STD_LOGIC;
		sclr	:	IN STD_LOGIC := '0';
		sload	:	IN STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
 BEGIN

	loop0 : FOR i IN 0 TO 4 GENERATE 
		wire_cntr2_w_lg_w_lg_sset334w335w(i) <= wire_cntr2_w_lg_sset334w(0) AND data(i);
	END GENERATE loop0;
	wire_cntr2_w_lg_clk_en342w(0) <= clk_en AND wire_cntr2_w_lg_w_lg_w_lg_cnt_en339w340w341w(0);
	loop2 : FOR i IN 0 TO 4 GENERATE 
		wire_cntr2_w_lg_sset336w(i) <= sset AND s_val(i);
	END GENERATE loop2;
	wire_cntr2_w_lg_external_cin332w(0) <= NOT external_cin;
	wire_cntr2_w_lg_sset334w(0) <= NOT sset;
	loop3 : FOR i IN 0 TO 4 GENERATE 
		wire_cntr2_w_lg_w_lg_sset336w337w(i) <= wire_cntr2_w_lg_sset336w(i) OR wire_cntr2_w_lg_w_lg_sset334w335w(i);
	END GENERATE loop3;
	wire_cntr2_w_lg_w_lg_w_lg_cnt_en339w340w341w(0) <= wire_cntr2_w_lg_w_lg_cnt_en339w340w(0) OR sload;
	wire_cntr2_w_lg_w_lg_cnt_en339w340w(0) <= wire_cntr2_w_lg_cnt_en339w(0) OR sset;
	wire_cntr2_w_lg_cnt_en339w(0) <= cnt_en OR sclr;
	wire_cntr2_w_lg_sset338w(0) <= sset OR sload;
	aclr_actual <= '0';
	clk_en <= '1';
	data <= (OTHERS => '0');
	external_cin <= '1';
	lsb_cin <= '0';
	q <= safe_q;
	s_val <= "11111";
	safe_q <= wire_counter_reg_bit20a_regout;
	sload <= '0';
	sset <= '0';
	updown_dir <= '1';
	updown_lsb <= updown_dir;
	updown_other_bits <= (wire_cntr2_w_lg_external_cin332w(0) OR updown_dir);
	counter_comb_bita_0 :  stratixii_lcell_comb
	  GENERIC MAP (
		EXTENDED_LUT => "OFF",
		LUT_MASK => "0000000000000000000000000000000000000000000000001010101010101010",
		SHARED_ARITH => "OFF"
	  )
	  PORT MAP ( 
		cin => lsb_cin,
		cout => wire_counter_comb_bita_0cout,
		dataa => wire_counter_reg_bit20a_regout(0),
		datab => updown_lsb,
		sumout => wire_counter_comb_bita_0sumout
	  );
	counter_comb_bita_1 :  stratixii_lcell_comb
	  GENERIC MAP (
		EXTENDED_LUT => "OFF",
		LUT_MASK => "0000000000000000010101010101010100000000000000000011001100110011",
		SHARED_ARITH => "OFF"
	  )
	  PORT MAP ( 
		cin => wire_counter_comb_bita_0cout,
		cout => wire_counter_comb_bita_1cout,
		dataa => wire_counter_reg_bit20a_regout(1),
		datab => updown_other_bits,
		sumout => wire_counter_comb_bita_1sumout
	  );
	counter_comb_bita_2 :  stratixii_lcell_comb
	  GENERIC MAP (
		EXTENDED_LUT => "OFF",
		LUT_MASK => "0000000000000000010101010101010100000000000000000011001100110011",
		SHARED_ARITH => "OFF"
	  )
	  PORT MAP ( 
		cin => wire_counter_comb_bita_1cout,
		cout => wire_counter_comb_bita_2cout,
		dataa => wire_counter_reg_bit20a_regout(2),
		datab => updown_other_bits,
		sumout => wire_counter_comb_bita_2sumout
	  );
	counter_comb_bita_3 :  stratixii_lcell_comb
	  GENERIC MAP (
		EXTENDED_LUT => "OFF",
		LUT_MASK => "0000000000000000010101010101010100000000000000000011001100110011",
		SHARED_ARITH => "OFF"
	  )
	  PORT MAP ( 
		cin => wire_counter_comb_bita_2cout,
		cout => wire_counter_comb_bita_3cout,
		dataa => wire_counter_reg_bit20a_regout(3),
		datab => updown_other_bits,
		sumout => wire_counter_comb_bita_3sumout
	  );
	counter_comb_bita_4 :  stratixii_lcell_comb
	  GENERIC MAP (
		EXTENDED_LUT => "OFF",
		LUT_MASK => "0000000000000000010101010101010100000000000000000011001100110011",
		SHARED_ARITH => "OFF"
	  )
	  PORT MAP ( 
		cin => wire_counter_comb_bita_3cout,
		dataa => wire_counter_reg_bit20a_regout(4),
		datab => updown_other_bits,
		sumout => wire_counter_comb_bita_4sumout
	  );
	wire_counter_reg_bit20a_adatasdata <= wire_cntr2_w_lg_w_lg_sset336w337w;
	loop8 : FOR i IN 0 TO 4 GENERATE
		wire_counter_reg_bit20a_ena(i) <= wire_cntr2_w_lg_clk_en342w(0);
	END GENERATE loop8;
	loop9 : FOR i IN 0 TO 4 GENERATE
		wire_counter_reg_bit20a_sload(i) <= wire_cntr2_w_lg_sset338w(0);
	END GENERATE loop9;
	counter_reg_bit20a_0 :  stratixii_lcell_ff
	  PORT MAP ( 
		aclr => aclr_actual,
		adatasdata => wire_counter_reg_bit20a_adatasdata(0),
		clk => clock,
		datain => wire_counter_comb_bita_0sumout,
		ena => wire_counter_reg_bit20a_ena(0),
		regout => wire_counter_reg_bit20a_regout(0),
		sclr => sclr,
		sload => wire_counter_reg_bit20a_sload(0)
	  );
	counter_reg_bit20a_1 :  stratixii_lcell_ff
	  PORT MAP ( 
		aclr => aclr_actual,
		adatasdata => wire_counter_reg_bit20a_adatasdata(1),
		clk => clock,
		datain => wire_counter_comb_bita_1sumout,
		ena => wire_counter_reg_bit20a_ena(1),
		regout => wire_counter_reg_bit20a_regout(1),
		sclr => sclr,
		sload => wire_counter_reg_bit20a_sload(1)
	  );
	counter_reg_bit20a_2 :  stratixii_lcell_ff
	  PORT MAP ( 
		aclr => aclr_actual,
		adatasdata => wire_counter_reg_bit20a_adatasdata(2),
		clk => clock,
		datain => wire_counter_comb_bita_2sumout,
		ena => wire_counter_reg_bit20a_ena(2),
		regout => wire_counter_reg_bit20a_regout(2),
		sclr => sclr,
		sload => wire_counter_reg_bit20a_sload(2)
	  );
	counter_reg_bit20a_3 :  stratixii_lcell_ff
	  PORT MAP ( 
		aclr => aclr_actual,
		adatasdata => wire_counter_reg_bit20a_adatasdata(3),
		clk => clock,
		datain => wire_counter_comb_bita_3sumout,
		ena => wire_counter_reg_bit20a_ena(3),
		regout => wire_counter_reg_bit20a_regout(3),
		sclr => sclr,
		sload => wire_counter_reg_bit20a_sload(3)
	  );
	counter_reg_bit20a_4 :  stratixii_lcell_ff
	  PORT MAP ( 
		aclr => aclr_actual,
		adatasdata => wire_counter_reg_bit20a_adatasdata(4),
		clk => clock,
		datain => wire_counter_comb_bita_4sumout,
		ena => wire_counter_reg_bit20a_ena(4),
		regout => wire_counter_reg_bit20a_regout(4),
		sclr => sclr,
		sload => wire_counter_reg_bit20a_sload(4)
	  );

 END RTL; --alt_remote_cntr_c88


--lpm_counter DEVICE_FAMILY="Stratix II" lpm_direction="UP" lpm_width=4 clock cnt_en q sclr
--VERSION_BEGIN 6.0 cbx_cycloneii 2006:02:07:15:19:20:SJ cbx_lpm_add_sub 2006:01:09:11:17:20:SJ cbx_lpm_compare 2006:01:09:11:15:40:SJ cbx_lpm_counter 2006:03:23:14:19:24:SJ cbx_lpm_decode 2006:01:09:11:16:44:SJ cbx_mgl 2006:05:17:10:06:16:SJ cbx_stratix 2006:05:17:09:28:32:SJ cbx_stratixii 2006:03:03:09:35:36:SJ  VERSION_END

 LIBRARY stratixii;
 USE stratixii.all;

--synthesis_resources = lut 4 reg 4 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  alt_remote_cntr_b88 IS 
	 PORT 
	 ( 
		 clock	:	IN  STD_LOGIC;
		 cnt_en	:	IN  STD_LOGIC := '1';
		 q	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 sclr	:	IN  STD_LOGIC := '0'
	 ); 
 END alt_remote_cntr_b88;

 ARCHITECTURE RTL OF alt_remote_cntr_b88 IS

	 ATTRIBUTE synthesis_clearbox : boolean;
	 ATTRIBUTE synthesis_clearbox OF RTL : ARCHITECTURE IS true;
	 SIGNAL  wire_counter_comb_bita_0cout	:	STD_LOGIC;
	 SIGNAL  wire_counter_comb_bita_1cout	:	STD_LOGIC;
	 SIGNAL  wire_counter_comb_bita_2cout	:	STD_LOGIC;
	 SIGNAL  wire_counter_comb_bita_0sumout	:	STD_LOGIC;
	 SIGNAL  wire_counter_comb_bita_1sumout	:	STD_LOGIC;
	 SIGNAL  wire_counter_comb_bita_2sumout	:	STD_LOGIC;
	 SIGNAL  wire_counter_comb_bita_3sumout	:	STD_LOGIC;
	 SIGNAL  wire_counter_reg_bit21a_adatasdata	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_counter_reg_bit21a_ena	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_counter_reg_bit21a_regout	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_counter_reg_bit21a_sload	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cntr3_w_lg_w_lg_sset345w346w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cntr3_w_lg_clk_en353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cntr3_w_lg_sset347w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cntr3_w_lg_external_cin343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cntr3_w_lg_sset345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cntr3_w_lg_w_lg_sset347w348w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cntr3_w_lg_w_lg_w_lg_cnt_en350w351w352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cntr3_w_lg_w_lg_cnt_en350w351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cntr3_w_lg_cnt_en350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_cntr3_w_lg_sset349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  aclr_actual :	STD_LOGIC;
	 SIGNAL  clk_en	:	STD_LOGIC;
	 SIGNAL  data	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  external_cin :	STD_LOGIC;
	 SIGNAL  lsb_cin :	STD_LOGIC;
	 SIGNAL  s_val :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  safe_q :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  sload	:	STD_LOGIC;
	 SIGNAL  sset	:	STD_LOGIC;
	 SIGNAL  updown_dir :	STD_LOGIC;
	 SIGNAL  updown_lsb :	STD_LOGIC;
	 SIGNAL  updown_other_bits :	STD_LOGIC;
	 COMPONENT  stratixii_lcell_comb
	 GENERIC 
	 (
		EXTENDED_LUT	:	STRING := "OFF";
		LUT_MASK	:	STD_LOGIC_VECTOR(63 DOWNTO 0);
		SHARED_ARITH	:	STRING := "OFF";
		lpm_type	:	STRING := "stratixii_lcell_comb"
	 );
	 PORT
	 ( 
		cin	:	IN STD_LOGIC := '0';
		combout	:	OUT STD_LOGIC;
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC := '0';
		datab	:	IN STD_LOGIC := '0';
		datac	:	IN STD_LOGIC := '0';
		datad	:	IN STD_LOGIC := '0';
		datae	:	IN STD_LOGIC := '0';
		dataf	:	IN STD_LOGIC := '0';
		datag	:	IN STD_LOGIC := '0';
		sharein	:	IN STD_LOGIC := '0';
		shareout	:	OUT STD_LOGIC;
		sumout	:	OUT STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  stratixii_lcell_ff
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		adatasdata	:	IN STD_LOGIC := '0';
		aload	:	IN STD_LOGIC := '0';
		clk	:	IN STD_LOGIC;
		datain	:	IN STD_LOGIC;
		ena	:	IN STD_LOGIC := '1';
		regout	:	OUT STD_LOGIC;
		sclr	:	IN STD_LOGIC := '0';
		sload	:	IN STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
 BEGIN

	loop10 : FOR i IN 0 TO 3 GENERATE 
		wire_cntr3_w_lg_w_lg_sset345w346w(i) <= wire_cntr3_w_lg_sset345w(0) AND data(i);
	END GENERATE loop10;
	wire_cntr3_w_lg_clk_en353w(0) <= clk_en AND wire_cntr3_w_lg_w_lg_w_lg_cnt_en350w351w352w(0);
	loop12 : FOR i IN 0 TO 3 GENERATE 
		wire_cntr3_w_lg_sset347w(i) <= sset AND s_val(i);
	END GENERATE loop12;
	wire_cntr3_w_lg_external_cin343w(0) <= NOT external_cin;
	wire_cntr3_w_lg_sset345w(0) <= NOT sset;
	loop13 : FOR i IN 0 TO 3 GENERATE 
		wire_cntr3_w_lg_w_lg_sset347w348w(i) <= wire_cntr3_w_lg_sset347w(i) OR wire_cntr3_w_lg_w_lg_sset345w346w(i);
	END GENERATE loop13;
	wire_cntr3_w_lg_w_lg_w_lg_cnt_en350w351w352w(0) <= wire_cntr3_w_lg_w_lg_cnt_en350w351w(0) OR sload;
	wire_cntr3_w_lg_w_lg_cnt_en350w351w(0) <= wire_cntr3_w_lg_cnt_en350w(0) OR sset;
	wire_cntr3_w_lg_cnt_en350w(0) <= cnt_en OR sclr;
	wire_cntr3_w_lg_sset349w(0) <= sset OR sload;
	aclr_actual <= '0';
	clk_en <= '1';
	data <= (OTHERS => '0');
	external_cin <= '1';
	lsb_cin <= '0';
	q <= safe_q;
	s_val <= "1111";
	safe_q <= wire_counter_reg_bit21a_regout;
	sload <= '0';
	sset <= '0';
	updown_dir <= '1';
	updown_lsb <= updown_dir;
	updown_other_bits <= (wire_cntr3_w_lg_external_cin343w(0) OR updown_dir);
	counter_comb_bita_0 :  stratixii_lcell_comb
	  GENERIC MAP (
		EXTENDED_LUT => "OFF",
		LUT_MASK => "0000000000000000000000000000000000000000000000001010101010101010",
		SHARED_ARITH => "OFF"
	  )
	  PORT MAP ( 
		cin => lsb_cin,
		cout => wire_counter_comb_bita_0cout,
		dataa => wire_counter_reg_bit21a_regout(0),
		datab => updown_lsb,
		sumout => wire_counter_comb_bita_0sumout
	  );
	counter_comb_bita_1 :  stratixii_lcell_comb
	  GENERIC MAP (
		EXTENDED_LUT => "OFF",
		LUT_MASK => "0000000000000000010101010101010100000000000000000011001100110011",
		SHARED_ARITH => "OFF"
	  )
	  PORT MAP ( 
		cin => wire_counter_comb_bita_0cout,
		cout => wire_counter_comb_bita_1cout,
		dataa => wire_counter_reg_bit21a_regout(1),
		datab => updown_other_bits,
		sumout => wire_counter_comb_bita_1sumout
	  );
	counter_comb_bita_2 :  stratixii_lcell_comb
	  GENERIC MAP (
		EXTENDED_LUT => "OFF",
		LUT_MASK => "0000000000000000010101010101010100000000000000000011001100110011",
		SHARED_ARITH => "OFF"
	  )
	  PORT MAP ( 
		cin => wire_counter_comb_bita_1cout,
		cout => wire_counter_comb_bita_2cout,
		dataa => wire_counter_reg_bit21a_regout(2),
		datab => updown_other_bits,
		sumout => wire_counter_comb_bita_2sumout
	  );
	counter_comb_bita_3 :  stratixii_lcell_comb
	  GENERIC MAP (
		EXTENDED_LUT => "OFF",
		LUT_MASK => "0000000000000000010101010101010100000000000000000011001100110011",
		SHARED_ARITH => "OFF"
	  )
	  PORT MAP ( 
		cin => wire_counter_comb_bita_2cout,
		dataa => wire_counter_reg_bit21a_regout(3),
		datab => updown_other_bits,
		sumout => wire_counter_comb_bita_3sumout
	  );
	wire_counter_reg_bit21a_adatasdata <= wire_cntr3_w_lg_w_lg_sset347w348w;
	loop18 : FOR i IN 0 TO 3 GENERATE
		wire_counter_reg_bit21a_ena(i) <= wire_cntr3_w_lg_clk_en353w(0);
	END GENERATE loop18;
	loop19 : FOR i IN 0 TO 3 GENERATE
		wire_counter_reg_bit21a_sload(i) <= wire_cntr3_w_lg_sset349w(0);
	END GENERATE loop19;
	counter_reg_bit21a_0 :  stratixii_lcell_ff
	  PORT MAP ( 
		aclr => aclr_actual,
		adatasdata => wire_counter_reg_bit21a_adatasdata(0),
		clk => clock,
		datain => wire_counter_comb_bita_0sumout,
		ena => wire_counter_reg_bit21a_ena(0),
		regout => wire_counter_reg_bit21a_regout(0),
		sclr => sclr,
		sload => wire_counter_reg_bit21a_sload(0)
	  );
	counter_reg_bit21a_1 :  stratixii_lcell_ff
	  PORT MAP ( 
		aclr => aclr_actual,
		adatasdata => wire_counter_reg_bit21a_adatasdata(1),
		clk => clock,
		datain => wire_counter_comb_bita_1sumout,
		ena => wire_counter_reg_bit21a_ena(1),
		regout => wire_counter_reg_bit21a_regout(1),
		sclr => sclr,
		sload => wire_counter_reg_bit21a_sload(1)
	  );
	counter_reg_bit21a_2 :  stratixii_lcell_ff
	  PORT MAP ( 
		aclr => aclr_actual,
		adatasdata => wire_counter_reg_bit21a_adatasdata(2),
		clk => clock,
		datain => wire_counter_comb_bita_2sumout,
		ena => wire_counter_reg_bit21a_ena(2),
		regout => wire_counter_reg_bit21a_regout(2),
		sclr => sclr,
		sload => wire_counter_reg_bit21a_sload(2)
	  );
	counter_reg_bit21a_3 :  stratixii_lcell_ff
	  PORT MAP ( 
		aclr => aclr_actual,
		adatasdata => wire_counter_reg_bit21a_adatasdata(3),
		clk => clock,
		datain => wire_counter_comb_bita_3sumout,
		ena => wire_counter_reg_bit21a_ena(3),
		regout => wire_counter_reg_bit21a_regout(3),
		sclr => sclr,
		sload => wire_counter_reg_bit21a_sload(3)
	  );

 END RTL; --alt_remote_cntr_b88

 LIBRARY stratixii;
 USE stratixii.all;

--synthesis_resources = lut 9 reg 38 stratixii_rublock 1 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  alt_remote_rmtupdt_srj IS 
	 PORT 
	 ( 
		 busy	:	OUT  STD_LOGIC;
		 clock	:	IN  STD_LOGIC;
		 data_out	:	OUT  STD_LOGIC_VECTOR (11 DOWNTO 0);
		 param	:	IN  STD_LOGIC_VECTOR (2 DOWNTO 0) := (OTHERS => '0');
		 pgmout	:	OUT  STD_LOGIC_VECTOR (2 DOWNTO 0);
		 read_param	:	IN  STD_LOGIC := '0';
		 reconfig	:	IN  STD_LOGIC := '0';
		 reset	:	IN  STD_LOGIC;
		 reset_timer	:	IN  STD_LOGIC := '0'
	 ); 
 END alt_remote_rmtupdt_srj;

 ARCHITECTURE RTL OF alt_remote_rmtupdt_srj IS

	 ATTRIBUTE synthesis_clearbox : boolean;
	 ATTRIBUTE synthesis_clearbox OF RTL : ARCHITECTURE IS true;
	 SIGNAL	 dffe10	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe11	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe12	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe13	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe14	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe15	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe16	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe17	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe18	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe19a	:	STD_LOGIC_VECTOR(2 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe4a	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := "000000000000"
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_dffe4a_CLRN	:	STD_LOGIC_VECTOR(11 DOWNTO 0);
	 SIGNAL	 wire_dffe4a_ENA	:	STD_LOGIC_VECTOR(11 DOWNTO 0);
	 SIGNAL	 dffe5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe6	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe7	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe8	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe9	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_cntr2_q	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_cntr3_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_sd1_pgmout	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_sd1_regout	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w215w218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w215w227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w221w222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_idle261w262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable53w58w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable53w94w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable53w98w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable53w62w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable53w66w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable53w70w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable53w74w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable53w78w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable53w82w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable53w86w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable53w90w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_load_enable53w54w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_idle261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_data274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_init_counter270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_post280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_pre_data269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rublock_regout_reg313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable59w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable99w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable55w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable63w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable67w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable71w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable75w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable79w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable83w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable87w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable91w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable95w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_data289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_init_counter286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_post_data295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_pre_data285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_param_decoder_param_latch_range211w229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_param_decoder_param_latch_range211w224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_shift_reg_clear50w51w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_bit_counter_all_done288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_bit_counter_param_start_match268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_clock303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_idle244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_data240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_init243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_init_counter242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_param260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_post239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_pre_data241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_select_shift_nloop312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable53w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_width_counter_all_done272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_width_counter_param_width_match273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_data235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_init238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_init_counter237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_load233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_param259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_post_data234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_pre_data236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_wait232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_param_decoder_param_latch_range211w212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_param_decoder_param_latch_range213w214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_param_decoder_param_latch_range216w217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_idle261w262w263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_clear50w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_reg_load_enable49w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  bit_counter_all_done :	STD_LOGIC;
	 SIGNAL  bit_counter_clear :	STD_LOGIC;
	 SIGNAL  bit_counter_enable :	STD_LOGIC;
	 SIGNAL  bit_counter_param_start :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  bit_counter_param_start_match :	STD_LOGIC;
	 SIGNAL  data_in	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  idle :	STD_LOGIC;
	 SIGNAL  param_decoder_param_latch :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  param_decoder_select :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  power_up :	STD_LOGIC;
	 SIGNAL  read_data :	STD_LOGIC;
	 SIGNAL  read_init :	STD_LOGIC;
	 SIGNAL  read_init_counter :	STD_LOGIC;
	 SIGNAL  read_post :	STD_LOGIC;
	 SIGNAL  read_pre_data :	STD_LOGIC;
	 SIGNAL  rublock_captnupdt :	STD_LOGIC;
	 SIGNAL  rublock_clock :	STD_LOGIC;
	 SIGNAL  rublock_reconfig :	STD_LOGIC;
	 SIGNAL  rublock_regin :	STD_LOGIC;
	 SIGNAL  rublock_regout :	STD_LOGIC;
	 SIGNAL  rublock_regout_reg :	STD_LOGIC;
	 SIGNAL  rublock_shiftnld :	STD_LOGIC;
	 SIGNAL  select_shift_nloop :	STD_LOGIC;
	 SIGNAL  shift_reg_clear :	STD_LOGIC;
	 SIGNAL  shift_reg_load_enable :	STD_LOGIC;
	 SIGNAL  shift_reg_serial_in :	STD_LOGIC;
	 SIGNAL  shift_reg_serial_out :	STD_LOGIC;
	 SIGNAL  shift_reg_shift_enable :	STD_LOGIC;
	 SIGNAL  start_bit_decoder_out :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  start_bit_decoder_param_select :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  w102w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w111w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w121w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w12w :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  w132w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w141w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w152w :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  w165w :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  w176w :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  w187w :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  w199w :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  w329w :	STD_LOGIC;
	 SIGNAL  w36w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  width_counter_all_done :	STD_LOGIC;
	 SIGNAL  width_counter_clear :	STD_LOGIC;
	 SIGNAL  width_counter_enable :	STD_LOGIC;
	 SIGNAL  width_counter_param_width :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  width_counter_param_width_match :	STD_LOGIC;
	 SIGNAL  width_decoder_out :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  width_decoder_param_select :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  write_data :	STD_LOGIC;
	 SIGNAL  write_init :	STD_LOGIC;
	 SIGNAL  write_init_counter :	STD_LOGIC;
	 SIGNAL  write_load :	STD_LOGIC;
	 SIGNAL  write_param	:	STD_LOGIC;
	 SIGNAL  write_post_data :	STD_LOGIC;
	 SIGNAL  write_pre_data :	STD_LOGIC;
	 SIGNAL  write_wait :	STD_LOGIC;
	 SIGNAL  wire_w_data_in_range57w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range97w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range52w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range61w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range65w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range69w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range73w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range77w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range81w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range85w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range89w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_data_in_range93w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_param_decoder_param_latch_range211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_param_decoder_param_latch_range213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_param_decoder_param_latch_range216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  alt_remote_cntr_c88
	 PORT
	 ( 
		clock	:	IN  STD_LOGIC;
		cnt_en	:	IN  STD_LOGIC := '1';
		q	:	OUT  STD_LOGIC_VECTOR(4 DOWNTO 0);
		sclr	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  alt_remote_cntr_b88
	 PORT
	 ( 
		clock	:	IN  STD_LOGIC;
		cnt_en	:	IN  STD_LOGIC := '1';
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		sclr	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  stratixii_rublock
	 GENERIC 
	 (
		operation_mode	:	STRING := "remote";
		sim_init_config	:	STRING := "factory";
		sim_init_page_select	:	NATURAL := 0;
		sim_init_status	:	NATURAL := 0;
		sim_init_watchdog_value	:	NATURAL := 0;
		lpm_type	:	STRING := "stratixii_rublock"
	 );
	 PORT
	 ( 
		captnupdt	:	IN STD_LOGIC;
		clk	:	IN STD_LOGIC;
		pgmout	:	OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
		rconfig	:	IN STD_LOGIC;
		regin	:	IN STD_LOGIC;
		regout	:	OUT STD_LOGIC;
		rsttimer	:	IN STD_LOGIC;
		shiftnld	:	IN STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	wire_w_lg_w215w218w(0) <= wire_w215w(0) AND wire_w_lg_w_param_decoder_param_latch_range216w217w(0);
	wire_w_lg_w215w227w(0) <= wire_w215w(0) AND wire_w_param_decoder_param_latch_range216w(0);
	wire_w_lg_w221w222w(0) <= wire_w221w(0) AND wire_w_lg_w_param_decoder_param_latch_range216w217w(0);
	wire_w_lg_w_lg_idle261w262w(0) <= wire_w_lg_idle261w(0) AND wire_w_lg_write_param259w(0);
	wire_w230w(0) <= wire_w_lg_w_param_decoder_param_latch_range211w229w(0) AND wire_w_param_decoder_param_latch_range216w(0);
	wire_w225w(0) <= wire_w_lg_w_param_decoder_param_latch_range211w224w(0) AND wire_w_lg_w_param_decoder_param_latch_range216w217w(0);
	wire_w_lg_w_lg_shift_reg_load_enable53w58w(0) <= wire_w_lg_shift_reg_load_enable53w(0) AND dffe4a(1);
	wire_w_lg_w_lg_shift_reg_load_enable53w94w(0) <= wire_w_lg_shift_reg_load_enable53w(0) AND dffe4a(10);
	wire_w_lg_w_lg_shift_reg_load_enable53w98w(0) <= wire_w_lg_shift_reg_load_enable53w(0) AND dffe4a(11);
	wire_w_lg_w_lg_shift_reg_load_enable53w62w(0) <= wire_w_lg_shift_reg_load_enable53w(0) AND dffe4a(2);
	wire_w_lg_w_lg_shift_reg_load_enable53w66w(0) <= wire_w_lg_shift_reg_load_enable53w(0) AND dffe4a(3);
	wire_w_lg_w_lg_shift_reg_load_enable53w70w(0) <= wire_w_lg_shift_reg_load_enable53w(0) AND dffe4a(4);
	wire_w_lg_w_lg_shift_reg_load_enable53w74w(0) <= wire_w_lg_shift_reg_load_enable53w(0) AND dffe4a(5);
	wire_w_lg_w_lg_shift_reg_load_enable53w78w(0) <= wire_w_lg_shift_reg_load_enable53w(0) AND dffe4a(6);
	wire_w_lg_w_lg_shift_reg_load_enable53w82w(0) <= wire_w_lg_shift_reg_load_enable53w(0) AND dffe4a(7);
	wire_w_lg_w_lg_shift_reg_load_enable53w86w(0) <= wire_w_lg_shift_reg_load_enable53w(0) AND dffe4a(8);
	wire_w_lg_w_lg_shift_reg_load_enable53w90w(0) <= wire_w_lg_shift_reg_load_enable53w(0) AND dffe4a(9);
	wire_w_lg_w_lg_shift_reg_load_enable53w54w(0) <= wire_w_lg_shift_reg_load_enable53w(0) AND shift_reg_serial_in;
	wire_w215w(0) <= wire_w_lg_w_param_decoder_param_latch_range211w212w(0) AND wire_w_lg_w_param_decoder_param_latch_range213w214w(0);
	wire_w221w(0) <= wire_w_lg_w_param_decoder_param_latch_range211w212w(0) AND wire_w_param_decoder_param_latch_range213w(0);
	wire_w_lg_idle261w(0) <= idle AND wire_w_lg_read_param260w(0);
	wire_w_lg_read_data274w(0) <= read_data AND wire_w_lg_width_counter_param_width_match273w(0);
	wire_w_lg_read_init_counter270w(0) <= read_init_counter AND wire_w_lg_bit_counter_param_start_match268w(0);
	wire_w_lg_read_post280w(0) <= read_post AND wire_w_lg_width_counter_all_done272w(0);
	wire_w_lg_read_pre_data269w(0) <= read_pre_data AND wire_w_lg_bit_counter_param_start_match268w(0);
	wire_w_lg_rublock_regout_reg313w(0) <= rublock_regout_reg AND wire_w_lg_select_shift_nloop312w(0);
	wire_w_lg_shift_reg_load_enable59w(0) <= shift_reg_load_enable AND wire_w_data_in_range57w(0);
	wire_w_lg_shift_reg_load_enable99w(0) <= shift_reg_load_enable AND wire_w_data_in_range97w(0);
	wire_w_lg_shift_reg_load_enable55w(0) <= shift_reg_load_enable AND wire_w_data_in_range52w(0);
	wire_w_lg_shift_reg_load_enable63w(0) <= shift_reg_load_enable AND wire_w_data_in_range61w(0);
	wire_w_lg_shift_reg_load_enable67w(0) <= shift_reg_load_enable AND wire_w_data_in_range65w(0);
	wire_w_lg_shift_reg_load_enable71w(0) <= shift_reg_load_enable AND wire_w_data_in_range69w(0);
	wire_w_lg_shift_reg_load_enable75w(0) <= shift_reg_load_enable AND wire_w_data_in_range73w(0);
	wire_w_lg_shift_reg_load_enable79w(0) <= shift_reg_load_enable AND wire_w_data_in_range77w(0);
	wire_w_lg_shift_reg_load_enable83w(0) <= shift_reg_load_enable AND wire_w_data_in_range81w(0);
	wire_w_lg_shift_reg_load_enable87w(0) <= shift_reg_load_enable AND wire_w_data_in_range85w(0);
	wire_w_lg_shift_reg_load_enable91w(0) <= shift_reg_load_enable AND wire_w_data_in_range89w(0);
	wire_w_lg_shift_reg_load_enable95w(0) <= shift_reg_load_enable AND wire_w_data_in_range93w(0);
	wire_w_lg_write_data289w(0) <= write_data AND wire_w_lg_width_counter_param_width_match273w(0);
	wire_w_lg_write_init_counter286w(0) <= write_init_counter AND wire_w_lg_bit_counter_param_start_match268w(0);
	wire_w_lg_write_post_data295w(0) <= write_post_data AND wire_w_lg_bit_counter_all_done288w(0);
	wire_w_lg_write_pre_data285w(0) <= write_pre_data AND wire_w_lg_bit_counter_param_start_match268w(0);
	wire_w_lg_w_param_decoder_param_latch_range211w229w(0) <= wire_w_param_decoder_param_latch_range211w(0) AND wire_w_lg_w_param_decoder_param_latch_range213w214w(0);
	wire_w_lg_w_param_decoder_param_latch_range211w224w(0) <= wire_w_param_decoder_param_latch_range211w(0) AND wire_w_param_decoder_param_latch_range213w(0);
	wire_w_lg_w_lg_shift_reg_clear50w51w(0) <= NOT wire_w_lg_shift_reg_clear50w(0);
	wire_w_lg_bit_counter_all_done288w(0) <= NOT bit_counter_all_done;
	wire_w_lg_bit_counter_param_start_match268w(0) <= NOT bit_counter_param_start_match;
	wire_w_lg_clock303w(0) <= NOT clock;
	wire_w_lg_idle244w(0) <= NOT idle;
	wire_w_lg_read_data240w(0) <= NOT read_data;
	wire_w_lg_read_init243w(0) <= NOT read_init;
	wire_w_lg_read_init_counter242w(0) <= NOT read_init_counter;
	wire_w_lg_read_param260w(0) <= NOT read_param;
	wire_w_lg_read_post239w(0) <= NOT read_post;
	wire_w_lg_read_pre_data241w(0) <= NOT read_pre_data;
	wire_w_lg_select_shift_nloop312w(0) <= NOT select_shift_nloop;
	wire_w_lg_shift_reg_load_enable53w(0) <= NOT shift_reg_load_enable;
	wire_w_lg_width_counter_all_done272w(0) <= NOT width_counter_all_done;
	wire_w_lg_width_counter_param_width_match273w(0) <= NOT width_counter_param_width_match;
	wire_w_lg_write_data235w(0) <= NOT write_data;
	wire_w_lg_write_init238w(0) <= NOT write_init;
	wire_w_lg_write_init_counter237w(0) <= NOT write_init_counter;
	wire_w_lg_write_load233w(0) <= NOT write_load;
	wire_w_lg_write_param259w(0) <= NOT write_param;
	wire_w_lg_write_post_data234w(0) <= NOT write_post_data;
	wire_w_lg_write_pre_data236w(0) <= NOT write_pre_data;
	wire_w_lg_write_wait232w(0) <= NOT write_wait;
	wire_w_lg_w_param_decoder_param_latch_range211w212w(0) <= NOT wire_w_param_decoder_param_latch_range211w(0);
	wire_w_lg_w_param_decoder_param_latch_range213w214w(0) <= NOT wire_w_param_decoder_param_latch_range213w(0);
	wire_w_lg_w_param_decoder_param_latch_range216w217w(0) <= NOT wire_w_param_decoder_param_latch_range216w(0);
	wire_w_lg_w_lg_w_lg_idle261w262w263w(0) <= wire_w_lg_w_lg_idle261w262w(0) OR write_wait;
	wire_w_lg_shift_reg_clear50w(0) <= shift_reg_clear OR reset;
	wire_w_lg_shift_reg_load_enable49w(0) <= shift_reg_load_enable OR shift_reg_shift_enable;
	bit_counter_all_done <= (((((NOT wire_cntr2_q(0)) AND wire_cntr2_q(1)) AND (NOT wire_cntr2_q(2))) AND wire_cntr2_q(3)) AND wire_cntr2_q(4));
	bit_counter_clear <= (read_init OR write_init);
	bit_counter_enable <= (((((((((read_init OR write_init) OR read_init_counter) OR write_init_counter) OR read_pre_data) OR write_pre_data) OR read_data) OR write_data) OR read_post) OR write_post_data);
	bit_counter_param_start <= start_bit_decoder_out;
	bit_counter_param_start_match <= (((((NOT w12w(0)) AND (NOT w12w(1))) AND (NOT w12w(2))) AND (NOT w12w(3))) AND (NOT w12w(4)));
	busy <= wire_w_lg_idle244w(0);
	data_in <= (OTHERS => '0');
	data_out <= dffe4a;
	idle <= dffe5;
	param_decoder_param_latch <= dffe19a;
	param_decoder_select <= ( wire_w230w & wire_w_lg_w215w227w & wire_w225w & wire_w_lg_w221w222w & wire_w_lg_w215w218w);
	pgmout <= wire_sd1_pgmout;
	power_up <= ((((((((((((wire_w_lg_idle244w(0) AND wire_w_lg_read_init243w(0)) AND wire_w_lg_read_init_counter242w(0)) AND wire_w_lg_read_pre_data241w(0)) AND wire_w_lg_read_data240w(0)) AND wire_w_lg_read_post239w(0)) AND wire_w_lg_write_init238w(0)) AND wire_w_lg_write_init_counter237w(0)) AND wire_w_lg_write_pre_data236w(0)) AND wire_w_lg_write_data235w(0)) AND wire_w_lg_write_post_data234w(0)) AND wire_w_lg_write_load233w(0)) AND wire_w_lg_write_wait232w(0));
	read_data <= dffe9;
	read_init <= dffe6;
	read_init_counter <= dffe7;
	read_post <= dffe10;
	read_pre_data <= dffe8;
	rublock_captnupdt <= wire_w_lg_write_load233w(0);
	rublock_clock <= ((wire_w_lg_clock303w(0) AND wire_w_lg_idle244w(0)) AND wire_w_lg_write_wait232w(0));
	rublock_reconfig <= (idle AND reconfig);
	rublock_regin <= (wire_w_lg_rublock_regout_reg313w(0) OR (shift_reg_serial_out AND select_shift_nloop));
	rublock_regout <= wire_sd1_regout;
	rublock_regout_reg <= dffe18;
	rublock_shiftnld <= (((((read_pre_data OR write_pre_data) OR read_data) OR write_data) OR read_post) OR write_post_data);
	select_shift_nloop <= (wire_w_lg_read_data274w(0) OR wire_w_lg_write_data289w(0));
	shift_reg_clear <= read_init;
	shift_reg_load_enable <= (idle AND write_param);
	shift_reg_serial_in <= (rublock_regout_reg AND select_shift_nloop);
	shift_reg_serial_out <= dffe4a(0);
	shift_reg_shift_enable <= (((read_data OR write_data) OR read_post) OR write_post_data);
	start_bit_decoder_out <= ((((w152w OR w165w) OR w176w) OR w187w) OR ( "0" & "0" & start_bit_decoder_param_select(4) & "0" & start_bit_decoder_param_select(4)));
	start_bit_decoder_param_select <= param_decoder_select;
	w102w <= ( "0" & width_decoder_param_select(0) & "0" & width_decoder_param_select(0));
	w111w <= ( width_decoder_param_select(1) & width_decoder_param_select(1) & "0" & "0");
	w121w <= ( "0" & "0" & "0" & width_decoder_param_select(2));
	w12w <= (wire_cntr2_q XOR bit_counter_param_start);
	w132w <= ( "0" & width_decoder_param_select(3) & width_decoder_param_select(3) & width_decoder_param_select(3));
	w141w <= ( "0" & "0" & "0" & width_decoder_param_select(4));
	w152w <= ( "0" & "0" & "0" & "0" & "0");
	w165w <= ( "0" & start_bit_decoder_param_select(1) & start_bit_decoder_param_select(1) & start_bit_decoder_param_select(1) & "0");
	w176w <= ( "0" & start_bit_decoder_param_select(2) & start_bit_decoder_param_select(2) & "0" & start_bit_decoder_param_select(2));
	w187w <= ( "0" & "0" & start_bit_decoder_param_select(3) & start_bit_decoder_param_select(3) & "0");
	w199w <= ( "0" & "0" & start_bit_decoder_param_select(4) & "0" & start_bit_decoder_param_select(4));
	w329w <= (idle AND (write_param OR read_param));
	w36w <= (wire_cntr3_q XOR width_counter_param_width);
	width_counter_all_done <= (((wire_cntr3_q(0) AND wire_cntr3_q(1)) AND (NOT wire_cntr3_q(2))) AND wire_cntr3_q(3));
	width_counter_clear <= (read_init OR write_init);
	width_counter_enable <= ((read_data OR write_data) OR read_post);
	width_counter_param_width <= width_decoder_out;
	width_counter_param_width_match <= ((((NOT w36w(0)) AND (NOT w36w(1))) AND (NOT w36w(2))) AND (NOT w36w(3)));
	width_decoder_out <= ((((w102w OR w111w) OR w121w) OR w132w) OR ( "0" & "0" & "0" & width_decoder_param_select(4)));
	width_decoder_param_select <= param_decoder_select;
	write_data <= dffe14;
	write_init <= dffe11;
	write_init_counter <= dffe12;
	write_load <= dffe16;
	write_param <= '0';
	write_post_data <= dffe15;
	write_pre_data <= dffe13;
	write_wait <= dffe17;
	wire_w_data_in_range57w(0) <= data_in(0);
	wire_w_data_in_range97w(0) <= data_in(10);
	wire_w_data_in_range52w(0) <= data_in(11);
	wire_w_data_in_range61w(0) <= data_in(1);
	wire_w_data_in_range65w(0) <= data_in(2);
	wire_w_data_in_range69w(0) <= data_in(3);
	wire_w_data_in_range73w(0) <= data_in(4);
	wire_w_data_in_range77w(0) <= data_in(5);
	wire_w_data_in_range81w(0) <= data_in(6);
	wire_w_data_in_range85w(0) <= data_in(7);
	wire_w_data_in_range89w(0) <= data_in(8);
	wire_w_data_in_range93w(0) <= data_in(9);
	wire_w_param_decoder_param_latch_range211w(0) <= param_decoder_param_latch(0);
	wire_w_param_decoder_param_latch_range213w(0) <= param_decoder_param_latch(1);
	wire_w_param_decoder_param_latch_range216w(0) <= param_decoder_param_latch(2);
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe10 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN dffe10 <= (((read_data AND width_counter_param_width_match) AND wire_w_lg_width_counter_all_done272w(0)) OR wire_w_lg_read_post280w(0));
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe11 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN dffe11 <= (idle AND write_param);
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe12 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN dffe12 <= write_init;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe13 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN dffe13 <= (wire_w_lg_write_init_counter286w(0) OR wire_w_lg_write_pre_data285w(0));
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe14 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN dffe14 <= (((write_init_counter AND bit_counter_param_start_match) OR (write_pre_data AND bit_counter_param_start_match)) OR (wire_w_lg_write_data289w(0) AND wire_w_lg_bit_counter_all_done288w(0)));
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe15 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN dffe15 <= (((write_data AND width_counter_param_width_match) AND wire_w_lg_bit_counter_all_done288w(0)) OR wire_w_lg_write_post_data295w(0));
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe16 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN dffe16 <= ((write_data AND bit_counter_all_done) OR (write_post_data AND bit_counter_all_done));
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe17 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN dffe17 <= write_load;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe18 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN dffe18 <= rublock_regout;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe19a <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (w329w = '1') THEN dffe19a <= param;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe4a_CLRN(0))
	BEGIN
		IF (wire_dffe4a_CLRN(0) = '0') THEN dffe4a(0) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ENA(0) = '1') THEN dffe4a(0) <= (wire_w_lg_shift_reg_load_enable59w(0) OR wire_w_lg_w_lg_shift_reg_load_enable53w58w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe4a_CLRN(1))
	BEGIN
		IF (wire_dffe4a_CLRN(1) = '0') THEN dffe4a(1) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ENA(1) = '1') THEN dffe4a(1) <= (wire_w_lg_shift_reg_load_enable63w(0) OR wire_w_lg_w_lg_shift_reg_load_enable53w62w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe4a_CLRN(2))
	BEGIN
		IF (wire_dffe4a_CLRN(2) = '0') THEN dffe4a(2) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ENA(2) = '1') THEN dffe4a(2) <= (wire_w_lg_shift_reg_load_enable67w(0) OR wire_w_lg_w_lg_shift_reg_load_enable53w66w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe4a_CLRN(3))
	BEGIN
		IF (wire_dffe4a_CLRN(3) = '0') THEN dffe4a(3) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ENA(3) = '1') THEN dffe4a(3) <= (wire_w_lg_shift_reg_load_enable71w(0) OR wire_w_lg_w_lg_shift_reg_load_enable53w70w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe4a_CLRN(4))
	BEGIN
		IF (wire_dffe4a_CLRN(4) = '0') THEN dffe4a(4) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ENA(4) = '1') THEN dffe4a(4) <= (wire_w_lg_shift_reg_load_enable75w(0) OR wire_w_lg_w_lg_shift_reg_load_enable53w74w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe4a_CLRN(5))
	BEGIN
		IF (wire_dffe4a_CLRN(5) = '0') THEN dffe4a(5) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ENA(5) = '1') THEN dffe4a(5) <= (wire_w_lg_shift_reg_load_enable79w(0) OR wire_w_lg_w_lg_shift_reg_load_enable53w78w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe4a_CLRN(6))
	BEGIN
		IF (wire_dffe4a_CLRN(6) = '0') THEN dffe4a(6) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ENA(6) = '1') THEN dffe4a(6) <= (wire_w_lg_shift_reg_load_enable83w(0) OR wire_w_lg_w_lg_shift_reg_load_enable53w82w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe4a_CLRN(7))
	BEGIN
		IF (wire_dffe4a_CLRN(7) = '0') THEN dffe4a(7) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ENA(7) = '1') THEN dffe4a(7) <= (wire_w_lg_shift_reg_load_enable87w(0) OR wire_w_lg_w_lg_shift_reg_load_enable53w86w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe4a_CLRN(8))
	BEGIN
		IF (wire_dffe4a_CLRN(8) = '0') THEN dffe4a(8) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ENA(8) = '1') THEN dffe4a(8) <= (wire_w_lg_shift_reg_load_enable91w(0) OR wire_w_lg_w_lg_shift_reg_load_enable53w90w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe4a_CLRN(9))
	BEGIN
		IF (wire_dffe4a_CLRN(9) = '0') THEN dffe4a(9) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ENA(9) = '1') THEN dffe4a(9) <= (wire_w_lg_shift_reg_load_enable95w(0) OR wire_w_lg_w_lg_shift_reg_load_enable53w94w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe4a_CLRN(10))
	BEGIN
		IF (wire_dffe4a_CLRN(10) = '0') THEN dffe4a(10) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ENA(10) = '1') THEN dffe4a(10) <= (wire_w_lg_shift_reg_load_enable99w(0) OR wire_w_lg_w_lg_shift_reg_load_enable53w98w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, wire_dffe4a_CLRN(11))
	BEGIN
		IF (wire_dffe4a_CLRN(11) = '0') THEN dffe4a(11) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (wire_dffe4a_ENA(11) = '1') THEN dffe4a(11) <= (wire_w_lg_shift_reg_load_enable55w(0) OR wire_w_lg_w_lg_shift_reg_load_enable53w54w(0));
			END IF;
		END IF;
	END PROCESS;
	loop71 : FOR i IN 0 TO 11 GENERATE
		wire_dffe4a_CLRN(i) <= wire_w_lg_w_lg_shift_reg_clear50w51w(0);
	END GENERATE loop71;
	loop72 : FOR i IN 0 TO 11 GENERATE
		wire_dffe4a_ENA(i) <= wire_w_lg_shift_reg_load_enable49w(0);
	END GENERATE loop72;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe5 <= '1';
		ELSIF (clock = '1' AND clock'event) THEN dffe5 <= (((wire_w_lg_w_lg_w_lg_idle261w262w263w(0) OR (read_data AND width_counter_all_done)) OR (read_post AND width_counter_all_done)) OR power_up);
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe6 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN dffe6 <= (idle AND read_param);
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe7 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN dffe7 <= read_init;
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe8 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN dffe8 <= (wire_w_lg_read_init_counter270w(0) OR wire_w_lg_read_pre_data269w(0));
		END IF;
	END PROCESS;
	PROCESS (clock, reset)
	BEGIN
		IF (reset = '1') THEN dffe9 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN dffe9 <= (((read_init_counter AND bit_counter_param_start_match) OR (read_pre_data AND bit_counter_param_start_match)) OR (wire_w_lg_read_data274w(0) AND wire_w_lg_width_counter_all_done272w(0)));
		END IF;
	END PROCESS;
	cntr2 :  alt_remote_cntr_c88
	  PORT MAP ( 
		clock => clock,
		cnt_en => bit_counter_enable,
		q => wire_cntr2_q,
		sclr => bit_counter_clear
	  );
	cntr3 :  alt_remote_cntr_b88
	  PORT MAP ( 
		clock => clock,
		cnt_en => width_counter_enable,
		q => wire_cntr3_q,
		sclr => width_counter_clear
	  );
	sd1 :  stratixii_rublock
	  GENERIC MAP (
		operation_mode => "local",
		sim_init_config => "application",
		sim_init_page_select => 1,
		sim_init_status => 15,
		sim_init_watchdog_value => 0
	  )
	  PORT MAP ( 
		captnupdt => rublock_captnupdt,
		clk => rublock_clock,
		pgmout => wire_sd1_pgmout,
		rconfig => rublock_reconfig,
		regin => rublock_regin,
		regout => wire_sd1_regout,
		rsttimer => reset_timer,
		shiftnld => rublock_shiftnld
	  );

 END RTL; --alt_remote_rmtupdt_srj
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY alt_remote IS
	PORT
	(
		clock		: IN STD_LOGIC ;
		param		: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		read_param		: IN STD_LOGIC ;
		reconfig		: IN STD_LOGIC ;
		reset		: IN STD_LOGIC ;
		reset_timer		: IN STD_LOGIC ;
		busy		: OUT STD_LOGIC ;
		data_out		: OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
		pgmout		: OUT STD_LOGIC_VECTOR (2 DOWNTO 0)
	);
END alt_remote;


ARCHITECTURE RTL OF alt_remote IS

	ATTRIBUTE synthesis_clearbox: boolean;
	ATTRIBUTE synthesis_clearbox OF RTL: ARCHITECTURE IS TRUE;
	SIGNAL sub_wire0	: STD_LOGIC ;
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (11 DOWNTO 0);
	SIGNAL sub_wire2	: STD_LOGIC_VECTOR (2 DOWNTO 0);



	COMPONENT alt_remote_rmtupdt_srj
	PORT (
			reconfig	: IN STD_LOGIC ;
			param	: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
			reset_timer	: IN STD_LOGIC ;
			read_param	: IN STD_LOGIC ;
			reset	: IN STD_LOGIC ;
			busy	: OUT STD_LOGIC ;
			clock	: IN STD_LOGIC ;
			data_out	: OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
			pgmout	: OUT STD_LOGIC_VECTOR (2 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	busy    <= sub_wire0;
	data_out    <= sub_wire1(11 DOWNTO 0);
	pgmout    <= sub_wire2(2 DOWNTO 0);

	alt_remote_rmtupdt_srj_component : alt_remote_rmtupdt_srj
	PORT MAP (
		reconfig => reconfig,
		param => param,
		reset_timer => reset_timer,
		read_param => read_param,
		reset => reset,
		clock => clock,
		busy => sub_wire0,
		data_out => sub_wire1,
		pgmout => sub_wire2
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix II"
-- Retrieval info: PRIVATE: SIM_INIT_CONFIG_COMBO STRING "APPLICATION"
-- Retrieval info: PRIVATE: SIM_INIT_PAGE_SELECT_COMBO STRING "1"
-- Retrieval info: PRIVATE: SIM_INIT_STAT_BIT0_CHECK STRING "1"
-- Retrieval info: PRIVATE: SIM_INIT_STAT_BIT1_CHECK STRING "1"
-- Retrieval info: PRIVATE: SIM_INIT_STAT_BIT2_CHECK STRING "1"
-- Retrieval info: PRIVATE: SIM_INIT_STAT_BIT3_CHECK STRING "1"
-- Retrieval info: PRIVATE: SIM_INIT_STAT_BIT4_CHECK STRING "0"
-- Retrieval info: PRIVATE: SIM_INIT_WATCHDOG_VALUE_EDIT STRING "1"
-- Retrieval info: PRIVATE: SUPPORT_WRITE_CHECK STRING "0"
-- Retrieval info: PRIVATE: WATCHDOG_ENABLE_CHECK STRING "0"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Stratix II"
-- Retrieval info: CONSTANT: OPERATION_MODE STRING "LOCAL"
-- Retrieval info: CONSTANT: SIM_INIT_CONFIG STRING "APPLICATION"
-- Retrieval info: CONSTANT: SIM_INIT_PAGE_SELECT NUMERIC "1"
-- Retrieval info: CONSTANT: SIM_INIT_STATUS NUMERIC "15"
-- Retrieval info: USED_PORT: busy 0 0 0 0 OUTPUT NODEFVAL "busy"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: USED_PORT: data_out 0 0 12 0 OUTPUT NODEFVAL "data_out[11..0]"
-- Retrieval info: USED_PORT: param 0 0 3 0 INPUT NODEFVAL "param[2..0]"
-- Retrieval info: USED_PORT: pgmout 0 0 3 0 OUTPUT NODEFVAL "pgmout[2..0]"
-- Retrieval info: USED_PORT: read_param 0 0 0 0 INPUT NODEFVAL "read_param"
-- Retrieval info: USED_PORT: reconfig 0 0 0 0 INPUT NODEFVAL "reconfig"
-- Retrieval info: USED_PORT: reset 0 0 0 0 INPUT NODEFVAL "reset"
-- Retrieval info: USED_PORT: reset_timer 0 0 0 0 INPUT NODEFVAL "reset_timer"
-- Retrieval info: CONNECT: @reset_timer 0 0 0 0 reset_timer 0 0 0 0
-- Retrieval info: CONNECT: @reset 0 0 0 0 reset 0 0 0 0
-- Retrieval info: CONNECT: @read_param 0 0 0 0 read_param 0 0 0 0
-- Retrieval info: CONNECT: pgmout 0 0 3 0 @pgmout 0 0 3 0
-- Retrieval info: CONNECT: data_out 0 0 12 0 @data_out 0 0 12 0
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: CONNECT: @param 0 0 3 0 param 0 0 3 0
-- Retrieval info: CONNECT: busy 0 0 0 0 @busy 0 0 0 0
-- Retrieval info: CONNECT: @reconfig 0 0 0 0 reconfig 0 0 0 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL alt_remote.vhd TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL alt_remote.inc TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL alt_remote.cmp FALSE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL alt_remote.bsf TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL alt_remote_inst.vhd FALSE FALSE
